module encoder_25x5(input logic[24:0] in
						 ,output logic[4:0] out);
	always_comb					 
		casez (in)		
			25'b0__0000_0000__0000_0000__0000_0001: out = 5'd24; 
			25'b0__0000_0000__0000_0000__0000_001?: out = 5'd23;  
			25'b0__0000_0000__0000_0000__0000_01??: out = 5'd22; 
			25'b0__0000_0000__0000_0000__0000_1???: out = 5'd21;  
			25'b0__0000_0000__0000_0000__0001_????: out = 5'd20;
			25'b0__0000_0000__0000_0000__001?_????: out = 5'd19;
			25'b0__0000_0000__0000_0000__01??_????: out = 5'd18; 
			25'b0__0000_0000__0000_0000__1???_????: out = 5'd17;
		
			25'b0__0000_0000__0000_0001__????_????: out = 5'd16;
			25'b0__0000_0000__0000_001?__????_????: out = 5'd15;
			25'b0__0000_0000__0000_01??__????_????: out = 5'd14;
			25'b0__0000_0000__0000_1???__????_????: out = 5'd13;
			25'b0__0000_0000__0001_????__????_????: out = 5'd12;		
			25'b0__0000_0000__001?_????__????_????: out = 5'd11;
			25'b0__0000_0000__01??_????__????_????: out = 5'd10;
			25'b0__0000_0000__1???_????__????_????: out = 5'd9;
			
			25'b0__0000_0001__????_????__????_????: out = 5'd8;
			25'b0__0000_001?__????_????__????_????: out = 5'd7;
			25'b0__0000_01??__????_????__????_????: out = 5'd6;
			25'b0__0000_1???__????_????__????_????: out = 5'd5;
			25'b0__0001_????__????_????__????_????: out = 5'd4;
			25'b0__001?_????__????_????__????_????: out = 5'd3;
			25'b0__01??_????__????_????__????_????: out = 5'd2;
			25'b0__1???_????__????_????__????_????: out = 5'd1;
			
			25'b1__????_????__????_????__????_????: out = 5'd0;
			default										  : out = 5'd31; 
		endcase
endmodule